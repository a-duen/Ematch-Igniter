CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 13 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
120 40 30 190 9
0 70 1025 733
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 70 1025 733
144179218 256
0
6 Title:
5 Name:
0
0
0
23
14 Opto Isolator~
173 502 164 0 4 9
0 3 7 6 8
0
0 0 880 782
7 OPTOISO
19 1 68 9
4 Cont
30 -9 58 -1
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 0
88 0 0 0 1 0 0 0
1 U
8953 0 0
0
0
7 Ground~
168 520 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 529 82 0 1 3
0 2
0
0 0 53344 512
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
9 Terminal~
194 430 126 0 1 3
0 3
0
0 0 49504 782
7 CONTpin
-26 -15 23 -7
2 T2
28 -17 42 -9
0
8 CONTpin;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6153 0 0
0
0
9 Terminal~
194 592 252 0 1 3
0 4
0
0 0 49504 270
7 readADC
-25 -15 24 -7
2 T3
-8 -25 6 -17
0
8 readADC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5394 0 0
0
0
9 Terminal~
194 189 207 0 1 3
0 5
0
0 0 49504 0
7 FIREpin
-24 -13 25 -5
2 T1
-7 -32 7 -24
0
8 FIREpin;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7734 0 0
0
0
10 Capacitor~
219 135 135 0 2 5
0 2 10
0
0 0 832 90
2 1u
14 0 28 8
7 Decoupl
11 -13 60 -5
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
2 +V
167 351 81 0 1 3
0 10
0
0 0 54240 0
3 11V
-10 -22 11 -14
7 BATTERY
-24 -32 25 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
7 Ground~
168 135 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
7 Ground~
168 387 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 324 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
7 Ground~
168 225 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 189 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
10 N-EMOS 3T~
219 378 243 0 3 7
0 6 9 2
0
0 0 832 0
5 BUZ11
13 1 48 9
6 MOSFET
11 -13 53 -5
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-220
7

0 2 3 1 2 3 1 0
77 0 0 256 1 1 0 0
1 Q
3363 0 0
0
0
14 Opto Isolator~
173 266 245 0 4 9
0 5 11 10 9
0
0 0 880 0
7 OPTOISO
-24 -28 25 -20
4 FIRE
-14 -38 14 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 0
88 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
9 Resistor~
219 592 108 0 4 5
0 7 2 0 -1
0
0 0 864 90
3 150
-26 -3 -5 5
7 optoRes
-52 -15 -3 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 484 99 0 4 5
0 3 2 0 -1
0
0 0 864 90
4 3.3k
4 -10 32 -2
7 pullRes
6 6 55 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 520 225 0 2 5
0 4 8
0
0 0 864 90
4 2.2k
8 0 36 8
5 divR1
13 -10 48 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 520 279 0 3 5
0 2 4 -1
0
0 0 864 90
3 470
5 0 26 8
5 divR2
14 -12 49 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 387 135 0 4 5
0 6 10 0 1
0
0 0 736 90
3 1.7
-24 -1 -3 7
6 EMATCH
-44 -15 -2 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 324 279 0 3 5
0 2 9 -1
0
0 0 864 90
4 2.2k
9 0 37 8
7 pullRes
4 -11 53 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 189 261 0 3 5
0 2 5 -1
0
0 0 864 90
4 3.3k
-35 11 -7 19
7 pullRes
-50 -1 -1 7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 225 279 0 3 5
0 2 11 -1
0
0 0 864 90
3 150
5 7 26 15
7 optoRes
6 -6 55 2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
24
3 0 6 0 0 4224 0 1 0 0 17 2
488 192
387 192
1 0 3 0 0 4224 0 4 0 0 3 2
440 125
484 125
1 1 3 0 0 0 0 17 1 0 0 3
484 117
484 138
488 138
1 0 2 0 0 4096 0 3 0 0 10 2
529 76
529 61
1 2 7 0 0 8320 0 16 1 0 0 3
592 126
592 138
512 138
4 2 8 0 0 8320 0 1 18 0 0 3
512 192
520 192
520 207
1 0 4 0 0 4224 0 5 0 0 9 2
580 251
520 251
1 1 2 0 0 0 0 2 19 0 0 2
520 309
520 297
1 2 4 0 0 0 0 18 19 0 0 2
520 243
520 261
2 2 2 0 0 8192 0 16 17 0 0 4
592 90
592 61
484 61
484 81
0 2 9 0 0 8320 0 0 14 12 0 3
324 257
324 252
360 252
4 2 9 0 0 0 0 15 21 0 0 3
292 257
324 257
324 261
1 0 5 0 0 4096 0 6 0 0 21 2
189 216
189 233
1 2 10 0 0 4096 0 8 20 0 0 3
351 90
387 90
387 117
1 3 10 0 0 12288 0 8 15 0 0 5
351 90
351 91
324 91
324 233
292 233
1 1 2 0 0 0 0 11 21 0 0 2
324 309
324 297
1 1 6 0 0 0 0 20 14 0 0 4
387 153
387 226
384 226
384 225
3 1 2 0 0 0 0 14 10 0 0 4
384 261
384 301
387 301
387 309
1 1 2 0 0 0 0 23 12 0 0 2
225 297
225 309
2 2 11 0 0 8320 0 23 15 0 0 3
225 261
225 257
238 257
1 2 5 0 0 4224 0 15 22 0 0 3
238 233
189 233
189 243
1 1 2 0 0 0 0 22 13 0 0 2
189 279
189 309
1 1 2 0 0 4224 0 7 9 0 0 2
135 144
135 309
2 0 10 0 0 8320 0 7 0 0 15 3
135 126
135 91
324 91
0
0
17 0 0
0
0
3 Vs1
0 3.3 3.3
0
0 0 0
3 0 1 4
0 4e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2951130 8419904 1357 101 0 0
77 66 647 246
688 71 1376 402
484 66
321 66
647 84
647 106
0 0
4.48037e-315 4.44803e-315 1.54261e-314 1.54703e-314 4.65474e-315 4.65474e-315
12409 0
4 5e-006 10
1
324 272
0 15 0 0 2	21 0 0 0
264620 1341504 100 100 0 0
0 0 0 0
21 143 182 213
0 0
0 0
0 66
0 66
0 0
0 0 0 0 0 0
12401 0
4 1 50
1
324 272
0 15 0 0 2	21 0 0 0
4395284 2259008 100 100 0 0
77 66 647 246
688 402 1376 733
647 66
77 66
647 66
647 246
0 0
0 0 0 0 0 0
12401 0
4 1 50
1
185 381
0 3 0 0 1	0 25 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
